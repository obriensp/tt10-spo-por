magic
tech sky130A
magscale 1 2
timestamp 1740960824
<< pwell >>
rect -2575 -2482 2575 2482
<< psubdiff >>
rect -2539 2412 -2443 2446
rect 2443 2412 2539 2446
rect -2539 2350 -2505 2412
rect 2505 2350 2539 2412
rect -2539 -2412 -2505 -2350
rect 2505 -2412 2539 -2350
rect -2539 -2446 -2443 -2412
rect 2443 -2446 2539 -2412
<< psubdiffcont >>
rect -2443 2412 2443 2446
rect -2539 -2350 -2505 2350
rect 2505 -2350 2539 2350
rect -2443 -2446 2443 -2412
<< xpolycontact >>
rect -2409 1884 -2271 2316
rect -2409 -2316 -2271 -1884
rect -2175 1884 -2037 2316
rect -2175 -2316 -2037 -1884
rect -1941 1884 -1803 2316
rect -1941 -2316 -1803 -1884
rect -1707 1884 -1569 2316
rect -1707 -2316 -1569 -1884
rect -1473 1884 -1335 2316
rect -1473 -2316 -1335 -1884
rect -1239 1884 -1101 2316
rect -1239 -2316 -1101 -1884
rect -1005 1884 -867 2316
rect -1005 -2316 -867 -1884
rect -771 1884 -633 2316
rect -771 -2316 -633 -1884
rect -537 1884 -399 2316
rect -537 -2316 -399 -1884
rect -303 1884 -165 2316
rect -303 -2316 -165 -1884
rect -69 1884 69 2316
rect -69 -2316 69 -1884
rect 165 1884 303 2316
rect 165 -2316 303 -1884
rect 399 1884 537 2316
rect 399 -2316 537 -1884
rect 633 1884 771 2316
rect 633 -2316 771 -1884
rect 867 1884 1005 2316
rect 867 -2316 1005 -1884
rect 1101 1884 1239 2316
rect 1101 -2316 1239 -1884
rect 1335 1884 1473 2316
rect 1335 -2316 1473 -1884
rect 1569 1884 1707 2316
rect 1569 -2316 1707 -1884
rect 1803 1884 1941 2316
rect 1803 -2316 1941 -1884
rect 2037 1884 2175 2316
rect 2037 -2316 2175 -1884
rect 2271 1884 2409 2316
rect 2271 -2316 2409 -1884
<< xpolyres >>
rect -2409 -1884 -2271 1884
rect -2175 -1884 -2037 1884
rect -1941 -1884 -1803 1884
rect -1707 -1884 -1569 1884
rect -1473 -1884 -1335 1884
rect -1239 -1884 -1101 1884
rect -1005 -1884 -867 1884
rect -771 -1884 -633 1884
rect -537 -1884 -399 1884
rect -303 -1884 -165 1884
rect -69 -1884 69 1884
rect 165 -1884 303 1884
rect 399 -1884 537 1884
rect 633 -1884 771 1884
rect 867 -1884 1005 1884
rect 1101 -1884 1239 1884
rect 1335 -1884 1473 1884
rect 1569 -1884 1707 1884
rect 1803 -1884 1941 1884
rect 2037 -1884 2175 1884
rect 2271 -1884 2409 1884
<< locali >>
rect -2539 2412 -2443 2446
rect 2443 2412 2539 2446
rect -2539 2350 -2505 2412
rect 2505 2350 2539 2412
rect -2539 -2412 -2505 -2350
rect 2505 -2412 2539 -2350
rect -2539 -2446 -2443 -2412
rect 2443 -2446 2539 -2412
<< viali >>
rect -2539 -1930 -2505 1930
rect 2505 -2171 2539 2171
rect -2255 -2446 2255 -2412
<< metal1 >>
rect 2499 2171 2545 2183
rect -2545 1930 -2499 1942
rect -2545 -1930 -2539 1930
rect -2505 -1930 -2499 1930
rect -2545 -1942 -2499 -1930
rect 2499 -2171 2505 2171
rect 2539 -2171 2545 2171
rect 2499 -2183 2545 -2171
rect -2267 -2412 2267 -2406
rect -2267 -2446 -2255 -2412
rect 2255 -2446 2267 -2412
rect -2267 -2452 2267 -2446
<< properties >>
string FIXED_BBOX -2522 -2429 2522 2429
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 19 m 1 nx 21 wmin 0.690 lmin 0.50 rho 2000 val 55.617k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 0 viagb 90 viagt 0 viagl 80 viagr 90
<< end >>
