magic
tech sky130A
magscale 1 2
timestamp 1740981720
<< locali >>
rect 74 7536 290 7770
rect 4490 7302 4706 7536
rect 74 7068 290 7302
rect 4490 6834 4706 7068
rect 74 6600 290 6834
rect 4490 6366 4706 6600
rect 74 6132 290 6366
rect 4490 5898 4706 6132
rect 74 5664 290 5898
rect 4490 5430 4706 5664
rect 74 5196 290 5430
rect 4490 4962 4706 5196
rect 74 4728 290 4962
rect 4490 4494 4706 4728
rect 74 4260 290 4494
rect 4490 4026 4706 4260
rect 74 3792 290 4026
rect 4490 3790 4706 3792
rect 4490 3558 4706 3574
rect 74 3324 290 3558
rect 4490 3090 4706 3324
<< viali >>
rect 4492 7702 4706 7840
rect 6044 5840 6080 5944
rect 5852 5702 5902 5754
rect 6044 5582 6080 5652
rect 4490 3574 4706 3790
rect 98 3010 290 3136
<< metal1 >>
rect -102 8106 -92 8406
rect 6460 8106 6470 8406
rect -92 3160 208 7976
rect -92 3136 314 3160
rect -92 3010 98 3136
rect 290 3010 314 3136
rect -92 2920 314 3010
rect -92 2898 208 2920
rect 508 2898 808 7976
rect 1108 2898 1408 7976
rect 1708 2898 2008 7976
rect 2308 2898 2608 7976
rect 2908 2898 3208 7976
rect 3508 2898 3808 7976
rect 4108 2898 4408 7976
rect 4480 7840 4718 8106
rect 4480 7702 4492 7840
rect 4706 7702 4718 7840
rect 4480 7690 4718 7702
rect 4908 4459 4918 8106
rect 5098 4959 5108 8106
rect 5308 5288 5318 8106
rect 5498 5288 5508 8106
rect 5708 6000 5718 8106
rect 5898 6086 5908 8106
rect 5898 6076 6456 6086
rect 6446 6000 6456 6076
rect 5708 5990 6456 6000
rect 6016 5944 6092 5960
rect 6016 5840 6044 5944
rect 6080 5840 6092 5944
rect 5840 5760 5914 5766
rect 5588 5754 5914 5760
rect 5588 5702 5852 5754
rect 5902 5702 5914 5754
rect 5588 5696 5914 5702
rect 5588 5404 5652 5696
rect 5840 5690 5914 5696
rect 6016 5760 6092 5840
rect 6016 5696 6180 5760
rect 6244 5696 6250 5760
rect 6016 5652 6092 5696
rect 6016 5582 6044 5652
rect 6080 5582 6092 5652
rect 6016 5574 6092 5582
rect 5728 5532 6460 5542
rect 5728 5456 5738 5532
rect 5728 5446 6270 5456
rect 6116 5404 6180 5410
rect 5588 5346 6116 5404
rect 5588 5340 6180 5346
rect 5308 5278 5508 5288
rect 5232 5046 5278 5052
rect 5390 5046 5436 5052
rect 5232 5000 5928 5046
rect 5166 4459 5176 4959
rect 5232 4418 5278 5000
rect 5310 4950 5356 5000
rect 5310 4418 5356 4506
rect 5390 4418 5436 5000
rect 5486 4459 5496 4959
rect 5828 4459 5838 4959
rect 5882 4418 5928 5000
rect 6116 4742 6180 4748
rect 5966 4684 6116 4742
rect 5966 4678 6180 4684
rect 5232 4388 5928 4418
rect 5208 4378 5928 4388
rect 5208 4372 5920 4378
rect 4478 3790 4712 3802
rect 4478 3574 4490 3790
rect 4706 3708 4712 3790
rect 5208 3762 5462 4372
rect 5310 3751 5356 3762
rect 4706 3662 5654 3708
rect 4706 3574 4712 3662
rect 4478 3562 4712 3574
rect -92 2756 4573 2898
rect 5082 2756 5582 3624
rect 6260 2756 6270 5446
rect 6450 2756 6460 5532
rect -102 2456 -92 2756
rect 6460 2456 6470 2756
<< via1 >>
rect -92 8106 6460 8406
rect 4918 4959 5098 8106
rect 5318 5288 5498 8106
rect 5718 6076 5898 8106
rect 5718 6000 6446 6076
rect 6180 5696 6244 5760
rect 5738 5456 6450 5532
rect 6116 5346 6180 5404
rect 4918 4459 5166 4959
rect 5496 4459 5828 4959
rect 6116 4684 6180 4742
rect 6270 2756 6450 5456
rect -92 2456 6460 2756
<< metal2 >>
rect -92 8406 6460 8416
rect -92 8096 4918 8106
rect 4908 4959 4918 8096
rect 5098 8096 5318 8106
rect 5098 5296 5108 8096
rect 5308 5296 5318 8096
rect 5098 5288 5318 5296
rect 5498 8096 5718 8106
rect 5498 5296 5508 8096
rect 5708 6000 5718 8096
rect 5898 8096 6460 8106
rect 5898 6086 5908 8096
rect 5898 6076 6456 6086
rect 6446 6000 6456 6076
rect 5708 5990 6456 6000
rect 6180 5760 6244 5766
rect 6306 5696 6315 5760
rect 6180 5690 6244 5696
rect 5728 5532 6460 5542
rect 5728 5456 5738 5532
rect 5728 5446 6270 5456
rect 6116 5405 6180 5414
rect 6110 5346 6116 5404
rect 6180 5346 6186 5404
rect 6116 5336 6180 5345
rect 5498 5288 5828 5296
rect 5098 5096 5828 5288
rect 5098 4959 5166 5096
rect 4918 4449 5166 4459
rect 5496 4959 5828 5096
rect 6116 4743 6180 4752
rect 6110 4684 6116 4742
rect 6180 4684 6186 4742
rect 6116 4674 6180 4683
rect 5496 4449 5828 4459
rect 6260 2766 6270 5446
rect -92 2756 6270 2766
rect 6450 2756 6460 5532
rect -92 2446 6460 2456
<< via2 >>
rect -92 8106 6460 8406
rect 6242 5696 6244 5760
rect 6244 5696 6306 5760
rect 6116 5404 6180 5405
rect 6116 5346 6180 5404
rect 6116 5345 6180 5346
rect 6116 4742 6180 4743
rect 6116 4684 6180 4742
rect 6116 4683 6180 4684
rect -92 2456 6460 2756
<< metal3 >>
rect -102 8406 6470 8411
rect -102 8106 -92 8406
rect 6460 8106 6470 8406
rect -102 8101 6470 8106
rect 6234 5760 6360 5768
rect 6234 5696 6242 5760
rect 6354 5696 6360 5760
rect 6234 5688 6360 5696
rect 6096 5410 6200 5424
rect 6096 5340 6111 5410
rect 6185 5340 6200 5410
rect 6096 5326 6200 5340
rect 6096 4748 6200 4762
rect 6096 4678 6111 4748
rect 6185 4678 6200 4748
rect 6096 4664 6200 4678
rect -92 2761 5988 2860
rect -102 2756 6470 2761
rect -102 2456 -92 2756
rect 6460 2456 6470 2756
rect -102 2451 6470 2456
<< via3 >>
rect -92 8106 6460 8406
rect 6290 5696 6306 5760
rect 6306 5696 6354 5760
rect 6111 5405 6185 5410
rect 6111 5345 6116 5405
rect 6116 5345 6180 5405
rect 6180 5345 6185 5405
rect 6111 5340 6185 5345
rect 6111 4743 6185 4748
rect 6111 4683 6116 4743
rect 6116 4683 6180 4743
rect 6180 4683 6185 4743
rect 6111 4678 6185 4683
rect -92 2456 6460 2756
<< metal4 >>
rect -93 8406 6461 8407
rect -93 8106 -92 8406
rect 6460 8106 6461 8406
rect -93 8105 6461 8106
rect 6289 5760 6355 5761
rect 6289 5696 6290 5760
rect 6354 5696 6355 5760
rect 6289 5695 6355 5696
rect 6290 5461 6354 5695
rect 6110 5410 6186 5411
rect 6110 5405 6111 5410
rect 5876 5345 6111 5405
rect 6110 5340 6111 5345
rect 6185 5340 6186 5410
rect 6270 5401 6470 5461
rect 6110 5339 6186 5340
rect 6110 4748 6186 4749
rect 6110 4743 6111 4748
rect 5896 4683 6111 4743
rect 6110 4678 6111 4683
rect 6185 4678 6186 4748
rect 6110 4677 6186 4678
rect -80 2757 5976 2874
rect -93 2756 6461 2757
rect -93 2456 -92 2756
rect 6460 2456 6461 2756
rect -93 2455 6461 2456
use sky130_fd_pr__cap_mim_m3_1_826CVA  sky130_fd_pr__cap_mim_m3_1_826CVA_0
timestamp 1740972924
transform 0 -1 2948 -1 0 5428
box -2571 -3040 2571 3040
use sky130_fd_sc_hd__tapvpwrvgnd_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6268 0 1 5494
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5824 0 1 5494
box -38 -48 406 592
use sky130_fd_pr__pfet_01v8_hvt_48T65H  XM1
timestamp 1740953238
transform 1 0 5904 0 1 4709
box -246 -469 246 469
use sky130_fd_pr__pfet_01v8_hvt_RUWLFK  XM5
timestamp 1740953238
transform 1 0 5333 0 1 4709
box -325 -469 325 469
use sky130_fd_pr__nfet_01v8_lvt_ZAB8C6  XM7
timestamp 1740957599
transform 0 -1 5332 1 0 3686
box -246 -460 246 460
use sky130_fd_pr__res_xhigh_po_0p69_JJJUAV  XR1
timestamp 1740960824
transform 0 1 2390 -1 0 5431
box -2575 -2482 2575 2482
<< labels >>
flabel metal4 -93 8105 6461 8407 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal4 -93 2455 6461 2757 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal4 6270 5401 6470 5461 0 FreeSans 256 0 0 0 reset_b
port 4 nsew
<< end >>
