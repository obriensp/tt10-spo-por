** sch_path: /home/sean/Development/HDL/tt10-spo-por/xschem/por.sch
.subckt por VDD VSS reset_b
*.PININFO VDD:I VSS:I reset_b:O
XC1 net1 VSS sky130_fd_pr__cap_mim_m3_1 W=18 L=42 m=1
x1 net1 VSS VSS VDD VDD net8 sky130_fd_sc_hd__inv_4
XR1 VSS net2 VSS sky130_fd_pr__res_xhigh_po_0p69 L=108 mult=1 m=1
XM5 net3 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=10 nf=4 m=1
XM6 net4 net4 net3 VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2.5 nf=1 m=1
XM7 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.5 W=2.5 nf=1 m=1
XR2 net2 VDD VSS sky130_fd_pr__res_xhigh_po_0p69 L=288 mult=1 m=1
XM1 net10 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2.5 nf=1 m=1
XM2 net5 net4 net10 VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2.5 nf=1 m=1
XM3 net5 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=0.5 W=10 nf=4 m=1
XM4 net6 net6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=5 nf=2 m=1
XM8 net7 net7 net6 VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2.5 nf=1 m=1
XM9 net7 net5 VSS VSS sky130_fd_pr__nfet_01v8 L=0.5 W=2.5 nf=1 m=1
XM10 net11 net6 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2.5 nf=1 m=1
XM11 net1 net7 net11 VDD sky130_fd_pr__pfet_01v8 L=0.5 W=2.5 nf=1 m=1
x2 net8 VSS VSS VDD VDD net9 sky130_fd_sc_hd__inv_1
x3 net9 VSS VSS VDD VDD net8 sky130_fd_sc_hd__inv_1
x4 net9 VSS VSS VDD VDD reset_b sky130_fd_sc_hd__buf_2
.ends
.end
