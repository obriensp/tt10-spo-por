magic
tech sky130A
magscale 1 2
timestamp 1740948629
<< pwell >>
rect -235 -34782 235 34782
<< psubdiff >>
rect -199 34712 -103 34746
rect 103 34712 199 34746
rect -199 34650 -165 34712
rect 165 34650 199 34712
rect -199 -34712 -165 -34650
rect 165 -34712 199 -34650
rect -199 -34746 -103 -34712
rect 103 -34746 199 -34712
<< psubdiffcont >>
rect -103 34712 103 34746
rect -199 -34650 -165 34650
rect 165 -34650 199 34650
rect -103 -34746 103 -34712
<< xpolycontact >>
rect -69 34184 69 34616
rect -69 -34616 69 -34184
<< xpolyres >>
rect -69 -34184 69 34184
<< locali >>
rect -199 34712 -103 34746
rect 103 34712 199 34746
rect -199 34650 -165 34712
rect 165 34650 199 34712
rect -199 -34712 -165 -34650
rect 165 -34712 199 -34650
rect -199 -34746 -103 -34712
rect 103 -34746 199 -34712
<< viali >>
rect -53 34201 53 34598
rect -53 -34598 53 -34201
<< metal1 >>
rect -59 34598 59 34610
rect -59 34201 -53 34598
rect 53 34201 59 34598
rect -59 34189 59 34201
rect -59 -34201 59 -34189
rect -59 -34598 -53 -34201
rect 53 -34598 59 -34201
rect -59 -34610 59 -34598
<< properties >>
string FIXED_BBOX -182 -34729 182 34729
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 342.0 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 991.849k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
