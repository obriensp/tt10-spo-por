magic
tech sky130A
timestamp 1740946518
<< checkpaint >>
rect -530 -130 1230 12282
<< metal4 >>
rect 100 500 300 11652
rect 400 500 600 11652
rect 3067 11052 3097 11152
rect 3343 11052 3373 11152
rect 3619 11052 3649 11152
rect 3895 11052 3925 11152
rect 4171 11052 4201 11152
rect 4447 11052 4477 11152
rect 4723 11052 4753 11152
rect 4999 11052 5029 11152
rect 5275 11052 5305 11152
rect 5551 11052 5581 11152
rect 5827 11052 5857 11152
rect 6103 11052 6133 11152
rect 6379 11052 6409 11152
rect 6655 11052 6685 11152
rect 6931 11052 6961 11152
rect 7207 11052 7237 11152
rect 7483 11052 7513 11152
rect 7759 11052 7789 11152
rect 8035 11052 8065 11152
rect 8311 11052 8341 11152
rect 8587 11052 8617 11152
rect 8863 11052 8893 11152
rect 9139 11052 9169 11152
rect 9415 11052 9445 11152
rect 9691 11052 9721 11152
rect 9967 11052 9997 11152
rect 10243 11052 10273 11152
rect 10519 11052 10549 11152
rect 10795 11052 10825 11152
rect 11071 11052 11101 11152
rect 11347 11052 11377 11152
rect 11623 11052 11653 11152
rect 11899 11052 11929 11152
rect 12175 11052 12205 11152
rect 12451 11052 12481 11152
rect 12727 11052 12757 11152
rect 13003 11052 13033 11152
rect 13279 11052 13309 11152
rect 13555 11052 13585 11152
rect 13831 11052 13861 11152
rect 14107 11052 14137 11152
rect 14383 11052 14413 11152
rect 14659 11052 14689 11152
<< labels >>
flabel metal4 s 14383 11052 14413 11152 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 11052 14689 11152 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 11052 14137 11152 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 13831 11052 13861 11152 0 FreeSans 240 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 13555 11052 13585 11152 0 FreeSans 240 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 13279 11052 13309 11152 0 FreeSans 240 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 13003 11052 13033 11152 0 FreeSans 240 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 12727 11052 12757 11152 0 FreeSans 240 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 12451 11052 12481 11152 0 FreeSans 240 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 12175 11052 12205 11152 0 FreeSans 240 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 11899 11052 11929 11152 0 FreeSans 240 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 11623 11052 11653 11152 0 FreeSans 240 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 11347 11052 11377 11152 0 FreeSans 240 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 11071 11052 11101 11152 0 FreeSans 240 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 10795 11052 10825 11152 0 FreeSans 240 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 10519 11052 10549 11152 0 FreeSans 240 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 10243 11052 10273 11152 0 FreeSans 240 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 9967 11052 9997 11152 0 FreeSans 240 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 9691 11052 9721 11152 0 FreeSans 240 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 4999 11052 5029 11152 0 FreeSans 240 90 0 0 uio_oe[0]
port 19 nsew signal output
flabel metal4 s 4723 11052 4753 11152 0 FreeSans 240 90 0 0 uio_oe[1]
port 20 nsew signal output
flabel metal4 s 4447 11052 4477 11152 0 FreeSans 240 90 0 0 uio_oe[2]
port 21 nsew signal output
flabel metal4 s 4171 11052 4201 11152 0 FreeSans 240 90 0 0 uio_oe[3]
port 22 nsew signal output
flabel metal4 s 3895 11052 3925 11152 0 FreeSans 240 90 0 0 uio_oe[4]
port 23 nsew signal output
flabel metal4 s 3619 11052 3649 11152 0 FreeSans 240 90 0 0 uio_oe[5]
port 24 nsew signal output
flabel metal4 s 3343 11052 3373 11152 0 FreeSans 240 90 0 0 uio_oe[6]
port 25 nsew signal output
flabel metal4 s 3067 11052 3097 11152 0 FreeSans 240 90 0 0 uio_oe[7]
port 26 nsew signal output
flabel metal4 s 7207 11052 7237 11152 0 FreeSans 240 90 0 0 uio_out[0]
port 27 nsew signal output
flabel metal4 s 6931 11052 6961 11152 0 FreeSans 240 90 0 0 uio_out[1]
port 28 nsew signal output
flabel metal4 s 6655 11052 6685 11152 0 FreeSans 240 90 0 0 uio_out[2]
port 29 nsew signal output
flabel metal4 s 6379 11052 6409 11152 0 FreeSans 240 90 0 0 uio_out[3]
port 30 nsew signal output
flabel metal4 s 6103 11052 6133 11152 0 FreeSans 240 90 0 0 uio_out[4]
port 31 nsew signal output
flabel metal4 s 5827 11052 5857 11152 0 FreeSans 240 90 0 0 uio_out[5]
port 32 nsew signal output
flabel metal4 s 5551 11052 5581 11152 0 FreeSans 240 90 0 0 uio_out[6]
port 33 nsew signal output
flabel metal4 s 5275 11052 5305 11152 0 FreeSans 240 90 0 0 uio_out[7]
port 34 nsew signal output
flabel metal4 s 9415 11052 9445 11152 0 FreeSans 240 90 0 0 uo_out[0]
port 35 nsew signal output
flabel metal4 s 9139 11052 9169 11152 0 FreeSans 240 90 0 0 uo_out[1]
port 36 nsew signal output
flabel metal4 s 8863 11052 8893 11152 0 FreeSans 240 90 0 0 uo_out[2]
port 37 nsew signal output
flabel metal4 s 8587 11052 8617 11152 0 FreeSans 240 90 0 0 uo_out[3]
port 38 nsew signal output
flabel metal4 s 8311 11052 8341 11152 0 FreeSans 240 90 0 0 uo_out[4]
port 39 nsew signal output
flabel metal4 s 8035 11052 8065 11152 0 FreeSans 240 90 0 0 uo_out[5]
port 40 nsew signal output
flabel metal4 s 7759 11052 7789 11152 0 FreeSans 240 90 0 0 uo_out[6]
port 41 nsew signal output
flabel metal4 s 7483 11052 7513 11152 0 FreeSans 240 90 0 0 uo_out[7]
port 42 nsew signal output
flabel metal4 100 500 300 11652 1 FreeSans 800 0 0 0 VDPWR
port 43 nsew power bidirectional
flabel metal4 400 500 600 11652 1 FreeSans 800 0 0 0 VGND
port 44 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 11152
<< end >>
