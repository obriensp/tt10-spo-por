magic
tech sky130A
magscale 1 2
timestamp 1740948629
<< pwell >>
rect -235 -6282 235 6282
<< psubdiff >>
rect -199 6212 -103 6246
rect 103 6212 199 6246
rect -199 6150 -165 6212
rect 165 6150 199 6212
rect -199 -6212 -165 -6150
rect 165 -6212 199 -6150
rect -199 -6246 -103 -6212
rect 103 -6246 199 -6212
<< psubdiffcont >>
rect -103 6212 103 6246
rect -199 -6150 -165 6150
rect 165 -6150 199 6150
rect -103 -6246 103 -6212
<< xpolycontact >>
rect -69 5684 69 6116
rect -69 -6116 69 -5684
<< xpolyres >>
rect -69 -5684 69 5684
<< locali >>
rect -199 6212 -103 6246
rect 103 6212 199 6246
rect -199 6150 -165 6212
rect 165 6150 199 6212
rect -199 -6212 -165 -6150
rect 165 -6212 199 -6150
rect -199 -6246 -103 -6212
rect 103 -6246 199 -6212
<< viali >>
rect -53 5701 53 6098
rect -53 -6098 53 -5701
<< metal1 >>
rect -59 6098 59 6110
rect -59 5701 -53 6098
rect 53 5701 59 6098
rect -59 5689 59 5701
rect -59 -5701 59 -5689
rect -59 -6098 -53 -5701
rect 53 -6098 59 -5701
rect -59 -6110 59 -6098
<< properties >>
string FIXED_BBOX -182 -6229 182 6229
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 57.0 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 165.762k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
