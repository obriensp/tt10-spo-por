magic
tech sky130A
magscale 1 2
timestamp 1740962336
<< locali >>
rect 74 7536 290 7770
rect 4490 7302 4706 7536
rect 74 7068 290 7302
rect 4490 6834 4706 7068
rect 74 6600 290 6834
rect 4490 6366 4706 6600
rect 74 6132 290 6366
rect 4490 5898 4706 6132
rect 74 5664 290 5898
rect 4490 5430 4706 5664
rect 74 5196 290 5430
rect 4490 4962 4706 5196
rect 74 4728 290 4962
rect 4490 4494 4706 4728
rect 74 4260 290 4494
rect 4490 4026 4706 4260
rect 74 3792 290 4026
rect 4490 3790 4706 3792
rect 4490 3558 4706 3574
rect 74 3324 290 3558
rect 4490 3090 4706 3324
<< viali >>
rect 4492 7702 4706 7840
rect 6036 5852 6070 5886
rect 5852 5714 5890 5750
rect 4490 3574 4706 3790
rect 98 3010 290 3136
<< metal1 >>
rect -632 8326 -432 8350
rect -102 8326 -92 8406
rect -632 8182 -92 8326
rect -632 8150 -432 8182
rect -102 8106 -92 8182
rect 6460 8331 6470 8406
rect 6636 8331 6802 8354
rect 6460 8211 6802 8331
rect 6460 8106 6470 8211
rect -92 3160 208 7976
rect -92 3136 314 3160
rect -92 3010 98 3136
rect 290 3010 314 3136
rect -92 2920 314 3010
rect -92 2898 208 2920
rect 508 2898 808 7976
rect 1108 2898 1408 7976
rect 1708 2898 2008 7976
rect 2308 2898 2608 7976
rect 2908 2898 3208 7976
rect 3508 2898 3808 7976
rect 4108 2898 4408 7976
rect 4480 7840 4718 8106
rect 4480 7702 4492 7840
rect 4706 7702 4718 7840
rect 4480 7690 4718 7702
rect 4908 4959 5108 8106
rect 5728 6066 6456 6086
rect 6636 6066 6802 8211
rect 7272 6534 7472 6624
rect 5728 6011 6802 6066
rect 5728 5990 6456 6011
rect 6636 6004 6802 6011
rect 7070 6494 7472 6534
rect 7070 5964 7110 6494
rect 7272 6424 7472 6494
rect 6512 5924 7110 5964
rect 6022 5890 6084 5898
rect 6512 5890 6552 5924
rect 6022 5886 6552 5890
rect 6022 5852 6036 5886
rect 6070 5852 6552 5886
rect 6022 5850 6552 5852
rect 6022 5838 6084 5850
rect 5840 5752 5902 5762
rect 6590 5752 6600 5852
rect 5840 5750 6600 5752
rect 5840 5714 5852 5750
rect 5890 5714 6600 5750
rect 5840 5712 6600 5714
rect 5840 5702 5902 5712
rect 6590 5612 6600 5712
rect 6840 5612 6850 5852
rect 5728 5521 6456 5542
rect 6612 5521 6772 5560
rect 5728 5467 6772 5521
rect 5728 5446 6456 5467
rect 5232 5046 5278 5052
rect 5390 5046 5436 5052
rect 5232 5000 5928 5046
rect 4908 4459 4918 4959
rect 5166 4459 5176 4959
rect 5232 4418 5278 5000
rect 5310 4950 5356 5000
rect 5310 4418 5356 4506
rect 5390 4418 5436 5000
rect 5486 4459 5496 4959
rect 5828 4459 5838 4959
rect 5882 4418 5928 5000
rect 6390 4748 6502 4760
rect 6390 4740 6401 4748
rect 5972 4666 6401 4740
rect 6390 4658 6401 4666
rect 6491 4658 6502 4748
rect 6390 4646 6502 4658
rect 5232 4388 5928 4418
rect 5208 4378 5928 4388
rect 5208 4372 5920 4378
rect 4478 3790 4712 3802
rect 4478 3574 4490 3790
rect 4706 3708 4712 3790
rect 5208 3762 5462 4372
rect 5310 3751 5356 3762
rect 4706 3662 5654 3708
rect 4706 3574 4712 3662
rect 4478 3562 4712 3574
rect -92 2756 4573 2898
rect 5082 2756 5582 3624
rect -728 2636 -528 2668
rect -102 2636 -92 2756
rect -728 2490 -92 2636
rect -728 2468 -528 2490
rect -102 2456 -92 2490
rect 6460 2653 6470 2756
rect 6612 2653 6772 5467
rect 6460 2535 6772 2653
rect 6460 2456 6470 2535
rect 6612 2512 6772 2535
<< via1 >>
rect -92 8106 6460 8406
rect 6600 5612 6840 5852
rect 4918 4459 5166 4959
rect 5496 4459 5828 4959
rect 6401 4658 6491 4748
rect -92 2456 6460 2756
<< metal2 >>
rect -92 8406 6460 8416
rect -92 8096 6460 8106
rect 6600 5852 6840 5862
rect 6600 5602 6840 5612
rect 4918 5096 5828 5296
rect 4918 4959 5166 5096
rect 4918 4449 5166 4459
rect 5496 4959 5828 5096
rect 6390 4748 6502 4760
rect 6390 4658 6401 4748
rect 6491 4658 6502 4748
rect 6390 4646 6502 4658
rect 5496 4449 5828 4459
rect -92 2756 6460 2766
rect -92 2446 6460 2456
<< via2 >>
rect -92 8106 6460 8406
rect 6600 5612 6840 5852
rect 6401 4658 6491 4748
rect -92 2456 6460 2756
<< metal3 >>
rect -102 8406 6470 8411
rect -102 8106 -92 8406
rect 6460 8106 6470 8406
rect -102 8101 6470 8106
rect 6590 5852 6850 5857
rect 6590 5612 6600 5852
rect 6840 5612 6850 5852
rect 6590 5607 6850 5612
rect 6390 4753 6502 4760
rect 6390 4653 6396 4753
rect 6496 4653 6502 4753
rect 6390 4646 6502 4653
rect -102 2756 6470 2761
rect -102 2456 -92 2756
rect 6460 2456 6470 2756
rect -102 2451 6470 2456
<< via3 >>
rect -92 8106 6460 8406
rect 6600 5612 6840 5852
rect 6396 4748 6496 4753
rect 6396 4658 6401 4748
rect 6401 4658 6491 4748
rect 6491 4658 6496 4748
rect 6396 4653 6496 4658
rect -92 2456 6460 2756
<< metal4 >>
rect -93 8406 6461 8407
rect -93 8106 -92 8406
rect 6460 8106 6461 8406
rect -93 8105 6461 8106
rect 6599 5852 6841 5853
rect 6599 5784 6600 5852
rect 6168 5686 6600 5784
rect 6599 5612 6600 5686
rect 6840 5612 6841 5852
rect 6599 5611 6841 5612
rect 6395 4753 6497 4754
rect 6395 4748 6396 4753
rect 6199 4658 6396 4748
rect 6395 4653 6396 4658
rect 6496 4653 6497 4753
rect 6395 4652 6497 4653
rect -88 2757 8 2876
rect -93 2756 6461 2757
rect -93 2456 -92 2756
rect 6460 2456 6461 2756
rect -93 2455 6461 2456
use sky130_fd_sc_hd__tapvpwrvgnd_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6268 0 1 5494
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5824 0 1 5494
box -38 -48 406 592
use sky130_fd_pr__cap_mim_m3_1_48F2XE  XC1
timestamp 1740948629
transform -1 0 3094 0 -1 5429
box -3186 -2571 3186 2571
use sky130_fd_pr__pfet_01v8_hvt_48T65H  XM1
timestamp 1740953238
transform 1 0 5904 0 1 4709
box -246 -469 246 469
use sky130_fd_pr__pfet_01v8_hvt_RUWLFK  XM5
timestamp 1740953238
transform 1 0 5333 0 1 4709
box -325 -469 325 469
use sky130_fd_pr__nfet_01v8_lvt_ZAB8C6  XM7
timestamp 1740957599
transform 0 -1 5332 1 0 3686
box -246 -460 246 460
use sky130_fd_pr__res_xhigh_po_0p69_JJJUAV  XR1
timestamp 1740960824
transform 0 1 2390 -1 0 5431
box -2575 -2482 2575 2482
<< labels >>
flabel metal1 -728 2468 -528 2668 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 -632 8150 -432 8350 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 7272 6424 7472 6624 0 FreeSans 256 0 0 0 reset_b
port 2 nsew
<< end >>
