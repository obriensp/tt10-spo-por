magic
tech sky130A
magscale 1 2
timestamp 1740948629
<< pwell >>
rect -2575 -2482 2575 2482
<< psubdiff >>
rect -2539 2412 -2443 2446
rect 2443 2412 2539 2446
rect -2539 2350 -2505 2412
rect 2505 2350 2539 2412
rect -2539 -2412 -2505 -2350
rect 2505 -2412 2539 -2350
rect -2539 -2446 -2443 -2412
rect 2443 -2446 2539 -2412
<< psubdiffcont >>
rect -2443 2412 2443 2446
rect -2539 -2350 -2505 2350
rect 2505 -2350 2539 2350
rect -2443 -2446 2443 -2412
<< xpolycontact >>
rect -2409 1884 -2271 2316
rect -2409 -2316 -2271 -1884
rect -2175 1884 -2037 2316
rect -2175 -2316 -2037 -1884
rect -1941 1884 -1803 2316
rect -1941 -2316 -1803 -1884
rect -1707 1884 -1569 2316
rect -1707 -2316 -1569 -1884
rect -1473 1884 -1335 2316
rect -1473 -2316 -1335 -1884
rect -1239 1884 -1101 2316
rect -1239 -2316 -1101 -1884
rect -1005 1884 -867 2316
rect -1005 -2316 -867 -1884
rect -771 1884 -633 2316
rect -771 -2316 -633 -1884
rect -537 1884 -399 2316
rect -537 -2316 -399 -1884
rect -303 1884 -165 2316
rect -303 -2316 -165 -1884
rect -69 1884 69 2316
rect -69 -2316 69 -1884
rect 165 1884 303 2316
rect 165 -2316 303 -1884
rect 399 1884 537 2316
rect 399 -2316 537 -1884
rect 633 1884 771 2316
rect 633 -2316 771 -1884
rect 867 1884 1005 2316
rect 867 -2316 1005 -1884
rect 1101 1884 1239 2316
rect 1101 -2316 1239 -1884
rect 1335 1884 1473 2316
rect 1335 -2316 1473 -1884
rect 1569 1884 1707 2316
rect 1569 -2316 1707 -1884
rect 1803 1884 1941 2316
rect 1803 -2316 1941 -1884
rect 2037 1884 2175 2316
rect 2037 -2316 2175 -1884
rect 2271 1884 2409 2316
rect 2271 -2316 2409 -1884
<< xpolyres >>
rect -2409 -1884 -2271 1884
rect -2175 -1884 -2037 1884
rect -1941 -1884 -1803 1884
rect -1707 -1884 -1569 1884
rect -1473 -1884 -1335 1884
rect -1239 -1884 -1101 1884
rect -1005 -1884 -867 1884
rect -771 -1884 -633 1884
rect -537 -1884 -399 1884
rect -303 -1884 -165 1884
rect -69 -1884 69 1884
rect 165 -1884 303 1884
rect 399 -1884 537 1884
rect 633 -1884 771 1884
rect 867 -1884 1005 1884
rect 1101 -1884 1239 1884
rect 1335 -1884 1473 1884
rect 1569 -1884 1707 1884
rect 1803 -1884 1941 1884
rect 2037 -1884 2175 1884
rect 2271 -1884 2409 1884
<< locali >>
rect -2539 2412 -2443 2446
rect 2443 2412 2539 2446
rect -2539 2350 -2505 2412
rect 2505 2350 2539 2412
rect -2539 -2412 -2505 -2350
rect 2505 -2412 2539 -2350
rect -2539 -2446 -2443 -2412
rect 2443 -2446 2539 -2412
<< viali >>
rect -2393 1901 -2287 2298
rect -2159 1901 -2053 2298
rect -1925 1901 -1819 2298
rect -1691 1901 -1585 2298
rect -1457 1901 -1351 2298
rect -1223 1901 -1117 2298
rect -989 1901 -883 2298
rect -755 1901 -649 2298
rect -521 1901 -415 2298
rect -287 1901 -181 2298
rect -53 1901 53 2298
rect 181 1901 287 2298
rect 415 1901 521 2298
rect 649 1901 755 2298
rect 883 1901 989 2298
rect 1117 1901 1223 2298
rect 1351 1901 1457 2298
rect 1585 1901 1691 2298
rect 1819 1901 1925 2298
rect 2053 1901 2159 2298
rect 2287 1901 2393 2298
rect -2393 -2298 -2287 -1901
rect -2159 -2298 -2053 -1901
rect -1925 -2298 -1819 -1901
rect -1691 -2298 -1585 -1901
rect -1457 -2298 -1351 -1901
rect -1223 -2298 -1117 -1901
rect -989 -2298 -883 -1901
rect -755 -2298 -649 -1901
rect -521 -2298 -415 -1901
rect -287 -2298 -181 -1901
rect -53 -2298 53 -1901
rect 181 -2298 287 -1901
rect 415 -2298 521 -1901
rect 649 -2298 755 -1901
rect 883 -2298 989 -1901
rect 1117 -2298 1223 -1901
rect 1351 -2298 1457 -1901
rect 1585 -2298 1691 -1901
rect 1819 -2298 1925 -1901
rect 2053 -2298 2159 -1901
rect 2287 -2298 2393 -1901
<< metal1 >>
rect -2399 2298 -2281 2310
rect -2399 1901 -2393 2298
rect -2287 1901 -2281 2298
rect -2399 1889 -2281 1901
rect -2165 2298 -2047 2310
rect -2165 1901 -2159 2298
rect -2053 1901 -2047 2298
rect -2165 1889 -2047 1901
rect -1931 2298 -1813 2310
rect -1931 1901 -1925 2298
rect -1819 1901 -1813 2298
rect -1931 1889 -1813 1901
rect -1697 2298 -1579 2310
rect -1697 1901 -1691 2298
rect -1585 1901 -1579 2298
rect -1697 1889 -1579 1901
rect -1463 2298 -1345 2310
rect -1463 1901 -1457 2298
rect -1351 1901 -1345 2298
rect -1463 1889 -1345 1901
rect -1229 2298 -1111 2310
rect -1229 1901 -1223 2298
rect -1117 1901 -1111 2298
rect -1229 1889 -1111 1901
rect -995 2298 -877 2310
rect -995 1901 -989 2298
rect -883 1901 -877 2298
rect -995 1889 -877 1901
rect -761 2298 -643 2310
rect -761 1901 -755 2298
rect -649 1901 -643 2298
rect -761 1889 -643 1901
rect -527 2298 -409 2310
rect -527 1901 -521 2298
rect -415 1901 -409 2298
rect -527 1889 -409 1901
rect -293 2298 -175 2310
rect -293 1901 -287 2298
rect -181 1901 -175 2298
rect -293 1889 -175 1901
rect -59 2298 59 2310
rect -59 1901 -53 2298
rect 53 1901 59 2298
rect -59 1889 59 1901
rect 175 2298 293 2310
rect 175 1901 181 2298
rect 287 1901 293 2298
rect 175 1889 293 1901
rect 409 2298 527 2310
rect 409 1901 415 2298
rect 521 1901 527 2298
rect 409 1889 527 1901
rect 643 2298 761 2310
rect 643 1901 649 2298
rect 755 1901 761 2298
rect 643 1889 761 1901
rect 877 2298 995 2310
rect 877 1901 883 2298
rect 989 1901 995 2298
rect 877 1889 995 1901
rect 1111 2298 1229 2310
rect 1111 1901 1117 2298
rect 1223 1901 1229 2298
rect 1111 1889 1229 1901
rect 1345 2298 1463 2310
rect 1345 1901 1351 2298
rect 1457 1901 1463 2298
rect 1345 1889 1463 1901
rect 1579 2298 1697 2310
rect 1579 1901 1585 2298
rect 1691 1901 1697 2298
rect 1579 1889 1697 1901
rect 1813 2298 1931 2310
rect 1813 1901 1819 2298
rect 1925 1901 1931 2298
rect 1813 1889 1931 1901
rect 2047 2298 2165 2310
rect 2047 1901 2053 2298
rect 2159 1901 2165 2298
rect 2047 1889 2165 1901
rect 2281 2298 2399 2310
rect 2281 1901 2287 2298
rect 2393 1901 2399 2298
rect 2281 1889 2399 1901
rect -2399 -1901 -2281 -1889
rect -2399 -2298 -2393 -1901
rect -2287 -2298 -2281 -1901
rect -2399 -2310 -2281 -2298
rect -2165 -1901 -2047 -1889
rect -2165 -2298 -2159 -1901
rect -2053 -2298 -2047 -1901
rect -2165 -2310 -2047 -2298
rect -1931 -1901 -1813 -1889
rect -1931 -2298 -1925 -1901
rect -1819 -2298 -1813 -1901
rect -1931 -2310 -1813 -2298
rect -1697 -1901 -1579 -1889
rect -1697 -2298 -1691 -1901
rect -1585 -2298 -1579 -1901
rect -1697 -2310 -1579 -2298
rect -1463 -1901 -1345 -1889
rect -1463 -2298 -1457 -1901
rect -1351 -2298 -1345 -1901
rect -1463 -2310 -1345 -2298
rect -1229 -1901 -1111 -1889
rect -1229 -2298 -1223 -1901
rect -1117 -2298 -1111 -1901
rect -1229 -2310 -1111 -2298
rect -995 -1901 -877 -1889
rect -995 -2298 -989 -1901
rect -883 -2298 -877 -1901
rect -995 -2310 -877 -2298
rect -761 -1901 -643 -1889
rect -761 -2298 -755 -1901
rect -649 -2298 -643 -1901
rect -761 -2310 -643 -2298
rect -527 -1901 -409 -1889
rect -527 -2298 -521 -1901
rect -415 -2298 -409 -1901
rect -527 -2310 -409 -2298
rect -293 -1901 -175 -1889
rect -293 -2298 -287 -1901
rect -181 -2298 -175 -1901
rect -293 -2310 -175 -2298
rect -59 -1901 59 -1889
rect -59 -2298 -53 -1901
rect 53 -2298 59 -1901
rect -59 -2310 59 -2298
rect 175 -1901 293 -1889
rect 175 -2298 181 -1901
rect 287 -2298 293 -1901
rect 175 -2310 293 -2298
rect 409 -1901 527 -1889
rect 409 -2298 415 -1901
rect 521 -2298 527 -1901
rect 409 -2310 527 -2298
rect 643 -1901 761 -1889
rect 643 -2298 649 -1901
rect 755 -2298 761 -1901
rect 643 -2310 761 -2298
rect 877 -1901 995 -1889
rect 877 -2298 883 -1901
rect 989 -2298 995 -1901
rect 877 -2310 995 -2298
rect 1111 -1901 1229 -1889
rect 1111 -2298 1117 -1901
rect 1223 -2298 1229 -1901
rect 1111 -2310 1229 -2298
rect 1345 -1901 1463 -1889
rect 1345 -2298 1351 -1901
rect 1457 -2298 1463 -1901
rect 1345 -2310 1463 -2298
rect 1579 -1901 1697 -1889
rect 1579 -2298 1585 -1901
rect 1691 -2298 1697 -1901
rect 1579 -2310 1697 -2298
rect 1813 -1901 1931 -1889
rect 1813 -2298 1819 -1901
rect 1925 -2298 1931 -1901
rect 1813 -2310 1931 -2298
rect 2047 -1901 2165 -1889
rect 2047 -2298 2053 -1901
rect 2159 -2298 2165 -1901
rect 2047 -2310 2165 -2298
rect 2281 -1901 2399 -1889
rect 2281 -2298 2287 -1901
rect 2393 -2298 2399 -1901
rect 2281 -2310 2399 -2298
<< properties >>
string FIXED_BBOX -2522 -2429 2522 2429
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 19 m 1 nx 21 wmin 0.690 lmin 0.50 rho 2000 val 55.617k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
