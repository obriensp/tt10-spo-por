magic
tech sky130A
magscale 1 2
timestamp 1740952864
<< pwell >>
rect -246 -460 246 460
<< nmoslvt >>
rect -50 -250 50 250
<< ndiff >>
rect -108 238 -50 250
rect -108 -238 -96 238
rect -62 -238 -50 238
rect -108 -250 -50 -238
rect 50 238 108 250
rect 50 -238 62 238
rect 96 -238 108 238
rect 50 -250 108 -238
<< ndiffc >>
rect -96 -238 -62 238
rect 62 -238 96 238
<< psubdiff >>
rect -210 390 -114 424
rect 114 390 210 424
rect -210 328 -176 390
rect 176 328 210 390
rect -210 -390 -176 -328
rect 176 -390 210 -328
rect -210 -424 -114 -390
rect 114 -424 210 -390
<< psubdiffcont >>
rect -114 390 114 424
rect -210 -328 -176 328
rect 176 -328 210 328
rect -114 -424 114 -390
<< poly >>
rect -50 322 50 338
rect -50 288 -34 322
rect 34 288 50 322
rect -50 250 50 288
rect -50 -288 50 -250
rect -50 -322 -34 -288
rect 34 -322 50 -288
rect -50 -338 50 -322
<< polycont >>
rect -34 288 34 322
rect -34 -322 34 -288
<< locali >>
rect -210 390 -114 424
rect 114 390 210 424
rect -210 351 -176 390
rect 176 328 210 390
rect -50 288 -34 322
rect 34 288 50 322
rect -96 238 -62 254
rect -96 -254 -62 -238
rect 62 238 96 254
rect 62 -254 96 -238
rect -50 -322 -34 -288
rect 34 -322 50 -288
rect -210 -390 -176 -351
rect 176 -390 210 -328
rect -210 -424 -114 -390
rect 114 -424 210 -390
<< viali >>
rect -210 328 -176 351
rect -210 -328 -176 328
rect -34 288 34 322
rect -96 -238 -62 238
rect 62 -238 96 238
rect -34 -322 34 -288
rect -210 -351 -176 -328
<< metal1 >>
rect -216 351 -170 363
rect -216 -351 -210 351
rect -176 -351 -170 351
rect -46 322 46 328
rect -46 288 -34 322
rect 34 288 46 322
rect -46 282 46 288
rect -102 238 -56 250
rect -102 -238 -96 238
rect -62 -238 -56 238
rect -102 -250 -56 -238
rect 56 238 102 250
rect 56 -238 62 238
rect 96 -238 102 238
rect 56 -250 102 -238
rect -46 -288 46 -282
rect -46 -322 -34 -288
rect 34 -322 46 -288
rect -46 -328 46 -322
rect -216 -363 -170 -351
<< properties >>
string FIXED_BBOX -193 -407 193 407
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 90 viagt 0
<< end >>
